`timescale 1ns / 1ps
module tx_top(
    input clk,                // Main clock input (drives the state machines)
    input rst,                // Reset input (active-high, resets the entire module)
    
    output tx_pin_out,        // Output signal that drives the transmission pin
    input [7:0] tx_data,      // 8-bit data to be transmitted
    input tx_buf_not_empty,   // Indicates if the TX buffer contains data to be sent
    output tx_read_buf        // Control signal to read data from the TX buffer
    );
    
    // Internal wires to connect the submodules
    wire tx_band_sig;         // Signal indicating when data transmission is active
    wire clk_bps;             // Baud rate clock signal, generated by tx_band_gen
    
    // Instance of the `tx_band_gen` module to generate the baud rate clock and transmission signal
    tx_band_gen tx_band_gen(
        .clk(clk),               // Connect main clock
        .rst(rst),               // Connect reset signal
        .band_sig(tx_band_sig),  // Transmission active signal
        .clk_bps(clk_bps)        // Baud rate clock signal
    );
    
    // Instance of the `tx_ctl` module to handle the transmission of the data
    tx_ctl tx_ctl(
        .clk(clk),               // Connect main clock
        .rst(rst),               // Connect reset signal
        .tx_clk_bps(clk_bps),    // Connect baud rate clock
        .tx_band_sig(tx_band_sig), // Transmission active signal
        .tx_pin_out(tx_pin_out), // The output pin for transmitting data
        .tx_data(tx_data),       // 8-bit data to be transmitted
        .tx_buf_not_empty(tx_buf_not_empty), // Signal indicating buffer has data
        .tx_read_buf(tx_read_buf)  // Control signal to read data from the buffer
    );
    
endmodule
